`ifndef _include_allocator_controller_
`define _include_allocator_controller_

/* Allocator Controller
 *
 * This module takes in image weights and filter weights and puts them in the
 * proper locations in memory for the DSP to process. These values must be
 * sent in order. This controller uses counters to track where in memory to
 * put the values, and whether there is enough space in memory for the values
 * to fit.
 *
 * The rule is that every image weight has a corresponding filter weight that
 * must be multiplied together, and that these will have the same counter
 * values. We'd like to store each weight in its own memory address, but we
 * don't have enough space for that, so everything is stored in 
 * (address % 512). The values that have been received are counted, and when
 * both issue and filter counters are at a value, the DSP is allowed to run
 * computations up to that value.
 *
 * As the DSP runs multiply/accumulates, it tracks the number of its own 
 * operations it has performed. Once the DSP has used a weight, we're allowed to
 * overwrite it with the next weight at (weight address + 512). So, as long as
 * the dsp counter is less than 512 behind the allocator counter, we can
 * continue accepting new data. As long as the allocator counter is ahead of
 * the DSP counter, we can continue DSP execution.
 *
 * This module handles the counters and memory writes for the "allocator" side
 * of the above process.
 */

/* TODO
 * 
 * 1. We need to write the appropriate stuff to result_ready and result_data
 * when the DSP has finished execution, which includes a few more operations
 * (add bias, leaky relu)
 *
 * 2. The control mechanism for blocking issue isn't currently implemented. We
 * need to track the counters and tell if we should stop issue based on those
 * numbers.
 */

module AllocatorController #(
        // Leaky relu for binary leak can be implemented quickly as a bitwise
        // shift. The leak factor has to be constant across all nets, so it's
        // here as a constant.
        // leak = 0: relu(x) = 0               | x<0, x | x>0
        // leak > 0: relu(x) = x[leak+17:leak] | x<0, x | x>0
        // Since it's a parameter, this won't generate a barrel shifter
        parameter filter_leak = 0
    )(
        // Data from issue stage. When X and Y are within the bounds of our
        // center +- filter halfsize, we'll accept the data
        input  wire [ 7:0] issue_a_x,
        input  wire [ 7:0] issue_a_y,
        input  wire [17:0] issue_a_data,
        input  wire        issue_a_blocked,
        
        // Here's our counter and the DSP's counter, as described above. The
        // block signal should be raised if we're far ahead of the DSP.
        output reg  [12:0] issue_a_alloc_counter,
        input  wire [12:0] issue_a_dsp_counter,
        output reg         issue_a_block,
        
        // Inputs of filter data, to come from _somewhere_.
        input  wire [17:0] filter_data,
        input  wire        filter_blocked,
        
        // Filter counter and filter dsp counter, as above. We don't generate
        // the filter issue counter, since it's the same for all allocators
        // and can be generated by the filter data source
        input  wire [12:0] filter_issue_counter,
        input  wire [12:0] filter_dsp_counter,
        output reg         filter_block,
        
        // Signals from the issue positioner describing which pixels we are
        // centered on. We should get a position signal before receiving any
        // data. When we do, center +- filter halfsize is our sensitive region.
        input  wire [ 7:0] center_x_input,
        input  wire [ 7:0] center_y_input,
        input  wire        center_write_enable,
        
        // Constant data about the filter, which we can use to compute the 
        // counter maximum and to apply the bias
        input  wire [ 2:0] filter_dim,
        input  wire [17:0] filter_bias,
        input  wire [12:0] filter_length,
        
        // RAMB write signals -- we need write access to the memory buffer
        output reg         ramb_a_write_en,
        output reg  [17:0] ramb_a_data,
        output reg  [ 9:0] ramb_a_addr,

        output reg         ramb_b_write_en,
        output reg  [17:0] ramb_b_data,
        output reg  [ 9:0] ramb_b_addr,
        
        // UNIMPLEMENTED but we should raise ready and set data once the DSP
        // is done with computation and we've run bias and relu
        // see TODO #1
        output reg         result_ready,
        output reg  [17:0] result_data,

        input  wire        clk,
        input  wire        rst
    );

    // Tracks the center of where this allocator is currently positioned
    // within the image
    // Note that the image is padded with zeroes of width filter_halfsize, so 
    // with an example 5x5 filter, the min of these values is (2, 2)
    reg [7:0] center_x;
    reg [7:0] center_y;

    // The halfsize of the filter -- distance of the edge of the filter from
    // the center, 2 for a 5x5 and 1 for a 3x3
    wire [1:0] filter_halfsize;
    assign filter_halfsize = (filter_dim == 3) ? 1 : 2;
    
    // Signals describing whether the current issue position is within our
    // range.
    wire issue_a_xrange;
    wire issue_a_yrange;
    wire issue_a_en;

    // issue_x is within range if it's within the bounds (center - halfsize,
    // center + halfsize)
    assign issue_a_xrange = (
        (issue_a_x >= center_x - filter_halfsize) &&
        (issue_a_x <= center_x + filter_halfsize)
    ) ? 1'b1 : 1'b0;
    // Same for y
    assign issue_a_yrange = (
        (issue_a_y >= center_y - filter_halfsize) &&
        (issue_a_y <= center_y + filter_halfsize)
    ) ? 1'b1 : 1'b0;
    
    // If we're in range of both X and Y, then the pixel is within our filter
    // bounds and we should read it into memory
    assign issue_a_en = (issue_a_xrange && issue_a_yrange);

    // Control the image data RAM writes and alloc counter
    always @(posedge clk) begin
        // Start off at 0, not blocking, and don't write anything to RAM
        if (rst) begin
            issue_a_alloc_counter <= 0;
            ramb_a_write_en <= 0;
            issue_a_block <= 0;

        // If the pixel is in range and not blocked / sitting still, we should 
        // accept it as our next value
        end else if (issue_a_en && !issue_a_blocked) begin
            // Here we need to check if issue_a_alloc_counter and 
            // issue_a_dsp_counter imply that we should block issue (i.e. if 
            // reading a new value into ramb would overwrite a value that the 
            // DSP hasn't been able to process yet
            // (same with filter)
            // see TODO #2
            
            // We're accepting the value as a memory write
            ramb_a_write_en <= 1;
            // Image data is mapped onto memory addresses [0-511]
            ramb_a_addr <= {1'b0, issue_a_alloc_counter[8:0]};
            // Read issue data into the memory write data line
            ramb_a_data <= issue_a_data;
            // And increment the counter to the next value
            issue_a_alloc_counter <= issue_a_alloc_counter + 1;
        
        // Otherwise, we're not accepting the data, turn off memory writes
        end else begin
            ramb_a_write_en <= 0;
        end
    end
    
    // Same as above block, except replace "image" with "filter"
    always @(posedge clk) begin
        // Initial: don't block, don't write anything
        if (rst) begin
            filter_block <= 0;
            ramb_b_write_en <= 0;

        // If filter isn't blocked, accept the data
        end else if (!filter_blocked) begin
            // See above and TODO #2
            
            // Write into memory
            ramb_b_write_en <= 1;
            // Filter is mapped to addresses [512-1023]
            ramb_b_addr <= {1'b1, filter_issue_counter[8:0]};
            // Set memory write data line
            ramb_b_data <= filter_data;
        
        // If we're blocked, turn off the memory writes
        end else begin
            ramb_b_write_en <= 0;
        end
    end

    // When the positioner raises our center_write_enable line, that's the
    // signal that we should accept the center_x and center_y signals
    // currently on the bus
    always @(posedge clk) begin
        if (center_write_enable) begin
            center_x <= center_x_input;
            center_y <= center_y_input;
        end
    end
    
    // This is a debug block (remove for synthesis)
    // It will make sure that certain module invariants aren't violated during
    // simulation
    always @(posedge clk) begin
        // center_x and center_y should be within the image bounds. The first
        // and last rows and columns are padding only
        if (center_x < filter_halfsize || center_x + filter_halfsize < center_x || 
            center_y < filter_halfsize || center_y + filter_halfsize < center_y) begin
            $display("Param error: Assigned an allocator to (%d, %d). Allowable range is (%d, %d) to (%d, %d).",
                center_x, center_y, filter_halfsize, filter_halfsize, -filter_halfsize, -filter_halfsize);
            $display("If you're sending an image, you need to pad it with 0's manually in the issue stage");
        end
    end
endmodule

 `endif // _include_allocator_controller_
