module ExecutorLane();

endmodule
