`ifndef _include_interface_
`define _include_interface_

/* Memory Interface
 *
 * This module is intended to expose the main image memory to the processing
 * unit / outside world. As you can see, there's nothing there. Maybe you can
 * write it!
 *
 * Xilinx seems to like using the AXI4 protocol to control this process. There
 * might be a tutorial online about how to make that happen.
 */

module Interface(

    );
`endif // _include_interface_
