module ExecutorDSP();
endmodule
