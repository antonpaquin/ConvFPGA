`ifndef _include_interface_
`define _include_interface_

module Interface(
    /*
    * This is intended to be the module that talks with the CPU to fill image
    * memroy. Do with it as you like.
    */

    );
`endif // _include_interface_
